;First Circuit LC:
V1  1  0  ac 1
R1	1  2  1000
R2  2  3  1000
L1  3  0  6.58mH
R3  2  0  1000
;.tran
.ac DEC 100  100  1000K
.probe
.end